`define REG_WIDTH 32
`define PRF_NUM_WIDTH 6
`define ARF_NUM_WIDTH 5
`define PRF_NUM 64
`define DEBUG
