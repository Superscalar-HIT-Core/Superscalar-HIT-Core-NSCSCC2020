`timescale 1ns / 1ps

module CP0(

    );
endmodule
