`timescale 1ns / 1ps

module IFU_test(

    );
endmodule
