`timescale 1ns / 1ps
`include "../defs.sv"
`include "../defines/defines.svh"
module TargetBuffer(
    input clk,
    input rst,
    input [31:0] br_PC,
    output [31:0] target_PC,
    input [79:0] ghist
);



endmodule