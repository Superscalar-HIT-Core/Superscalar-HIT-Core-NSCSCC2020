`timescale 1ns / 1ps
`include "defines/defines.svh"
module exception(

    );
endmodule
