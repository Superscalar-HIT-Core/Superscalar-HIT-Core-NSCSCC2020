`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2020/07/19 23:05:36
// Design Name: 
// Module Name: MDU
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
`include "defines/defines.svh"

module MDU(
    input UOPBundle uopHi,
    input UOPBundle uopLo,

    output PRFwInfo wbData,
    FU_ROB.fu   mdu_rob
);

    

endmodule
