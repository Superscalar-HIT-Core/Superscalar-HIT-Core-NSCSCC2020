`timescale 1ns / 1ps
`include "defines/defines.svh"
module pipeline(
    input clk,
    input rst
    );



endmodule
